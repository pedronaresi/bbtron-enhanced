module instructionMemory (addy, clock, RAMOuput, reset);
  input [9:0] addy;
  input clock;
  input reset;

  output [31:0] RAMOuput;

  integer firstClock = 0;

  reg [31:0] instructionRAM [150:0];

  always @ (addy or reset) begin
    if (reset) begin
      // Algoritmmo a ser executado pelo processador
		
		instructionRAM[0] = 32'b010111_00000000000000000001010010; 	// Jump to Main
		instructionRAM[1] = 32'b001011_00011_00011_0000000000000111; 	// addi
		instructionRAM[2] = 32'b100000_00111_01011_0000000000000000; 	// mov
		instructionRAM[3] = 32'b100000_01000_01100_0000000000000000; 	// mov
		instructionRAM[4] = 32'b100000_01001_01101_0000000000000000; 	// mov
		instructionRAM[5] = 32'b010000_00011_01100_0000000000000000; 	// sw
		instructionRAM[6] = 32'b000000_01011_01100_10101_00000000000; 	// add
		instructionRAM[7] = 32'b001111_10101_10101_0000000000000000; 	// lw
		instructionRAM[8] = 32'b010000_00011_10101_1111111111111111; 	// sw
		instructionRAM[9] = 32'b001011_01100_10110_0000000000000001; 	// addi
		instructionRAM[10] = 32'b010000_00011_10110_1111111111111110; 	// sw
		instructionRAM[11] = 32'b001111_00011_01110_1111111111111110; 	// lw
		instructionRAM[12] = 32'b011100_01110_01101_0000000000011000; 	// blt
		instructionRAM[13] = 32'b000000_01011_01110_10111_00000000000; 	// add
		instructionRAM[14] = 32'b001111_10111_10111_0000000000000000; 	// lw
		instructionRAM[15] = 32'b001111_00011_01111_1111111111111111; 	// lw
		instructionRAM[16] = 32'b011100_10111_01111_0000000000010101; 	// blt
		instructionRAM[17] = 32'b000000_01011_01110_11000_00000000000; 	// add
		instructionRAM[18] = 32'b001111_11000_11000_0000000000000000; 	// lw
		instructionRAM[19] = 32'b010000_00011_11000_1111111111111111; 	// sw
		instructionRAM[20] = 32'b010000_00011_01110_0000000000000000; 	// sw
		instructionRAM[21] = 32'b001011_01110_11001_0000000000000001; 	// addi
		instructionRAM[22] = 32'b010000_00011_11001_1111111111111110; 	// sw
		instructionRAM[23] = 32'b010111_00000000000000000000001011; 	// j
		instructionRAM[24] = 32'b001111_00011_10000_0000000000000000; 	// lw
		instructionRAM[25] = 32'b100000_10000_00001_0000000000000000; 	// mov
		instructionRAM[26] = 32'b011011_00000_11111_0000000000000000; 	// jr
		instructionRAM[27] = 32'b001011_00011_00011_0000000000000111; 	// addi
		instructionRAM[28] = 32'b100000_00111_01011_0000000000000000; 	// mov
		instructionRAM[29] = 32'b100000_01000_01100_0000000000000000; 	// mov
		instructionRAM[30] = 32'b100000_01001_01101_0000000000000000; 	// mov
		instructionRAM[31] = 32'b010000_00011_01100_1111111111111110; 	// sw
		instructionRAM[32] = 32'b001100_01101_10101_0000000000000001; 	// subi
		instructionRAM[33] = 32'b001111_00011_01110_1111111111111110; 	// lw
		instructionRAM[34] = 32'b011100_01110_10101_0000000000111011; 	// blt
		instructionRAM[35] = 32'b010001_00011_00100_1111111111111011; 	// la
		instructionRAM[36] = 32'b100000_01110_01000_0000000000000000; 	// mov
		instructionRAM[37] = 32'b100000_01101_01001_0000000000000000; 	// mov
		instructionRAM[38] = 32'b010000_00011_11111_0000000000000001; 	// sw
		instructionRAM[39] = 32'b011010_00000000000000000000000001; 	// jal
		instructionRAM[40] = 32'b001100_00011_00011_0000000000000111; 	// subi
		instructionRAM[41] = 32'b001111_00011_11111_0000000000000001; 	// lw
		instructionRAM[42] = 32'b100000_00001_10110_0000000000000000; 	// mov
		instructionRAM[43] = 32'b010000_00011_10110_1111111111111111; 	// sw
		instructionRAM[44] = 32'b001111_00011_01111_1111111111111111; 	// lw
		instructionRAM[45] = 32'b000000_01011_01111_10111_00000000000; 	// add
		instructionRAM[46] = 32'b001111_10111_10111_0000000000000000; 	// lw
		instructionRAM[47] = 32'b010000_00011_10111_0000000000000000; 	// sw
		instructionRAM[48] = 32'b001111_00011_10000_1111111111111110; 	// lw
		instructionRAM[49] = 32'b000000_01011_10000_11000_00000000000; 	// add
		instructionRAM[50] = 32'b001111_11000_11000_0000000000000000; 	// lw
		instructionRAM[51] = 32'b000000_01011_01111_11001_00000000000; 	// add
		instructionRAM[52] = 32'b010000_11001_11000_0000000000000000; 	// sw
		instructionRAM[53] = 32'b000000_01011_10000_11010_00000000000; 	// add
		instructionRAM[54] = 32'b001111_00011_10001_0000000000000000; 	// lw
		instructionRAM[55] = 32'b010000_11010_10001_0000000000000000; 	// sw
		instructionRAM[56] = 32'b001011_10000_11011_0000000000000001; 	// addi
		instructionRAM[57] = 32'b010000_00011_11011_1111111111111110; 	// sw
		instructionRAM[58] = 32'b010111_00000000000000000000100000; 	// j
		instructionRAM[59] = 32'b011011_00000_11111_0000000000000000; 	// jr
		instructionRAM[60] = 32'b001011_00011_00011_0000000000000011; 	// addi
		instructionRAM[61] = 32'b100000_00111_01011_0000000000000000; 	// mov
		instructionRAM[62] = 32'b100000_01000_01100_0000000000000000; 	// mov
		instructionRAM[63] = 32'b100001_00000_10101_0000000000000000; 	// li
		instructionRAM[64] = 32'b001001_01100_10101_0000000001000100; 	// beq
		instructionRAM[65] = 32'b100000_01011_00001_0000000000000000; 	// mov
		instructionRAM[66] = 32'b011011_00000_11111_0000000000000000; 	// jr
		instructionRAM[67] = 32'b010111_00000000000000000001010001; 	// j
		instructionRAM[68] = 32'b100000_01100_00111_0000000000000000; 	// mov
		instructionRAM[69] = 32'b001111_00011_01101_0000000000000000; 	// lw
		instructionRAM[70] = 32'b000111_01011_01101_10110_00000000000; 	// div
		instructionRAM[71] = 32'b000110_10110_01101_10111_00000000000; 	// mul
		instructionRAM[72] = 32'b000001_01011_10111_11000_00000000000; 	// sub
		instructionRAM[73] = 32'b100000_11000_01000_0000000000000000; 	// mov
		instructionRAM[74] = 32'b010000_00011_11111_0000000000000001; 	// sw
		instructionRAM[75] = 32'b011010_00000000000000000000111100; 	// jal
		instructionRAM[76] = 32'b001100_00011_00011_0000000000000011; 	// subi
		instructionRAM[77] = 32'b001111_00011_11111_0000000000000001; 	// lw
		instructionRAM[78] = 32'b100000_00001_11001_0000000000000000; 	// mov
		instructionRAM[79] = 32'b100000_11001_00001_0000000000000000; 	// mov
		instructionRAM[80] = 32'b011011_00000_11111_0000000000000000; 	// jr
		instructionRAM[81] = 32'b011011_00000_11111_0000000000000000; 	// jr
		instructionRAM[82] = 32'b001011_00011_00011_0000000000001101; 	// addi
		instructionRAM[83] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[84] = 32'b111111_00000_10101_0000000000000000; 	// in
		instructionRAM[85] = 32'b010000_00011_10101_1111111111111101; 	// sw
		instructionRAM[86] = 32'b001111_00011_01011_1111111111111101; 	// lw
		instructionRAM[87] = 32'b100001_00000_10110_0000000000000000; 	// li
		instructionRAM[88] = 32'b011110_01011_10110_0000000010010000; 	// bgt
		instructionRAM[89] = 32'b100001_00000_10111_0000000000000001; 	// li
		instructionRAM[90] = 32'b001001_01011_10111_0000000001111011; 	// beq
		instructionRAM[91] = 32'b100001_00000_11000_0000000000000000; 	// li
		instructionRAM[92] = 32'b010000_00011_11000_1111111111111110; 	// sw
		instructionRAM[93] = 32'b001111_00011_01100_1111111111111110; 	// lw
		instructionRAM[94] = 32'b100001_00000_11001_0000000000001010; 	// li
		instructionRAM[95] = 32'b011100_01100_11001_0000000001101000; 	// blt
		instructionRAM[96] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[97] = 32'b111111_00000_11010_0000000000000000; 	// in
		instructionRAM[98] = 32'b010001_00101_01101_0000000000000000; 	// la
		instructionRAM[99] = 32'b000000_01101_01100_11011_00000000000; 	// add
		instructionRAM[100] = 32'b010000_11011_11010_0000000000000000; 	// sw
		instructionRAM[101] = 32'b001011_01100_11100_0000000000000001; 	// addi
		instructionRAM[102] = 32'b010000_00011_11100_1111111111111110; 	// sw
		instructionRAM[103] = 32'b010111_00000000000000000001011101; 	// j
		instructionRAM[104] = 32'b010001_00011_01010_1111111111111101; 	// la
		instructionRAM[105] = 32'b100001_00000_01000_0000000000000000; 	// li
		instructionRAM[106] = 32'b100001_00000_01001_0000000000001010; 	// li
		instructionRAM[107] = 32'b011010_00000000000000000000011011; 	// jal
		instructionRAM[108] = 32'b100000_00001_11101_0000000000000000; 	// mov
		instructionRAM[109] = 32'b001100_00011_00011_0000000000000111; 	// subi
		instructionRAM[110] = 32'b100001_00000_11110_0000000000000000; 	// li
		instructionRAM[111] = 32'b010000_00011_11110_1111111111111110; 	// sw
		instructionRAM[112] = 32'b001111_00011_01110_1111111111111110; 	// lw
		instructionRAM[113] = 32'b100001_00000_10101_0000000000001010; 	// li
		instructionRAM[114] = 32'b011100_01110_10101_0000000001111010; 	// blt
		instructionRAM[115] = 32'b000000_01101_01110_10101_00000000000; 	// add
		instructionRAM[116] = 32'b001111_10101_10101_0000000000000000; 	// lw
		instructionRAM[117] = 32'b100000_10101_00111_0000000000000000; 	// mov
		instructionRAM[118] = 32'b111110_00000_00111_0000000000000000; 	// out
		instructionRAM[119] = 32'b001011_01110_10110_0000000000000001; 	// addi
		instructionRAM[120] = 32'b010000_00011_10110_1111111111111110; 	// sw
		instructionRAM[121] = 32'b010111_00000000000000000001110000; 	// j
		instructionRAM[122] = 32'b010111_00000000000000000010001100; 	// j
		instructionRAM[123] = 32'b100001_00000_10111_0000000000000010; 	// li
		instructionRAM[124] = 32'b001001_01011_10111_0000000010001100; 	// beq
		instructionRAM[125] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[126] = 32'b111111_00000_11000_0000000000000000; 	// in
		instructionRAM[127] = 32'b010000_00011_11000_1111111111111111; 	// sw
		instructionRAM[128] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[129] = 32'b111111_00000_11001_0000000000000000; 	// in
		instructionRAM[130] = 32'b010000_00011_11001_0000000000000000; 	// sw
		instructionRAM[131] = 32'b001111_00011_01111_1111111111111111; 	// lw
		instructionRAM[132] = 32'b100000_01111_00111_0000000000000000; 	// mov
		instructionRAM[133] = 32'b001111_00011_10000_0000000000000000; 	// lw
		instructionRAM[134] = 32'b100000_10000_01000_0000000000000000; 	// mov
		instructionRAM[135] = 32'b011010_00000000000000000000111100; 	// jal
		instructionRAM[136] = 32'b100000_00001_11010_0000000000000000; 	// mov
		instructionRAM[137] = 32'b001100_00011_00011_0000000000000011; 	// subi
		instructionRAM[138] = 32'b100000_11010_00111_0000000000000000; 	// mov
		instructionRAM[139] = 32'b111110_00000_00111_0000000000000000; 	// out
		instructionRAM[140] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[141] = 32'b111111_00000_11011_0000000000000000; 	// in
		instructionRAM[142] = 32'b010000_00011_11011_1111111111111101; 	// sw
		instructionRAM[143] = 32'b010111_00000000000000000001010110; 	// j
		instructionRAM[144] = 32'b011101_00000000000000000000000000; 	// halt
		
		/*instructionRAM[0] = 32'b010111_00000000000000000000000001; 	// Jump to Main
		instructionRAM[1] = 32'b001011_00011_00011_0000000000000000; 	// addi
		instructionRAM[2] = 32'b011101_00000000000000000000000000; 	// halt
		instructionRAM[3] = 32'b010101_00000_10101_0000000000000000; 	// in
		instructionRAM[4] = 32'b010000_00011_10101_0000000000000000; 	// sw
		instructionRAM[5] = 32'b001111_00011_01011_0000000000000000; 	// lw
		instructionRAM[6] = 32'b100000_01011_00111_0000000000000000; 	// mov
		instructionRAM[7] = 32'b010110_00111_000000000000000000000; 	// out
		instructionRAM[8] = 32'b011101_00000000000000000000000000; 	// halt*/

		
		/*
		instructionRAM[0] = 32'b010110_00000_000000000000000000000; //out R[0]
		instructionRAM[1] = 32'b010101_00000_00010_0000000000000000; //in R[2] <- X
		instructionRAM[2] = 32'b010110_00010_000000000000000000000;	//out R[2]
		instructionRAM[3] = 32'b010101_00000_00001_0000000000000000; //in R[1] <- 0
		instructionRAM[4] = 32'b010110_00001_000000000000000000000; //out R[1]
		instructionRAM[5] = 32'b010101_00000_00011_0000000000000000; //in R[3] <- 2
		instructionRAM[6] = 32'b010110_00011_000000000000000000000; //out R[3]
		instructionRAM[7] = 32'b010101_00000_00110_0000000000000000; //in R[6] <- 5
		instructionRAM[8] = 32'b010110_00110_000000000000000000000; //out R[6]
		
		instructionRAM[9] = 32'b010000_00000_00010_0000000000000001; //sw do R[2] no MEM[1]
		
		instructionRAM[10] = 32'b001001_00001_00110_0000000000010000; // beq R[1] e R[6]
		instructionRAM[11] = 32'b001101_00000_00010_0000000000000000; //inc R[2]
		instructionRAM[12] = 32'b000110_00011_00010_00010_00000000000; //mul R[2] = R[2] * R[3]
		instructionRAM[13] = 32'b010110_00010_000000000000000000000; //out R[2]
		instructionRAM[14] = 32'b001101_00000_00001_0000000000000000; //inc R[1]
		instructionRAM[15] = 32'b010111_00000000000000000000001010; //j INS[10]
		instructionRAM[16] = 32'b001111_00000_00100_0000000000000001; //lw do MEM[1] no R[4]
		
		instructionRAM[17] = 32'b000001_00100_00010_00101_00000000000; //sub R[5] = R[4] - R[2]
		instructionRAM[18] = 32'b010110_00101_000000000000000000000; //out R[5]
		instructionRAM[19] = 32'b011000_00101_000000000000000000000; // hlt
		*/
    end
  end

  assign RAMOuput = (instructionRAM[addy]);

endmodule // Memória de instrução
